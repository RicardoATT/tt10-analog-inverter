magic
tech sky130A
magscale 1 2
timestamp 1740547666
<< nwell >>
rect -241 -354 241 354
<< pmos >>
rect -45 -135 45 135
<< pdiff >>
rect -103 123 -45 135
rect -103 -123 -91 123
rect -57 -123 -45 123
rect -103 -135 -45 -123
rect 45 123 103 135
rect 45 -123 57 123
rect 91 -123 103 123
rect 45 -135 103 -123
<< pdiffc >>
rect -91 -123 -57 123
rect 57 -123 91 123
<< nsubdiff >>
rect -205 284 -109 318
rect 109 284 205 318
rect -205 222 -171 284
rect 171 222 205 284
rect -205 -284 -171 -222
rect 171 -284 205 -222
rect -205 -318 -109 -284
rect 109 -318 205 -284
<< nsubdiffcont >>
rect -109 284 109 318
rect -205 -222 -171 222
rect 171 -222 205 222
rect -109 -318 109 -284
<< poly >>
rect -45 216 45 232
rect -45 182 -29 216
rect 29 182 45 216
rect -45 135 45 182
rect -45 -182 45 -135
rect -45 -216 -29 -182
rect 29 -216 45 -182
rect -45 -232 45 -216
<< polycont >>
rect -29 182 29 216
rect -29 -216 29 -182
<< locali >>
rect -205 284 -109 318
rect 109 284 205 318
rect -205 222 -171 284
rect 171 222 205 284
rect -45 182 -29 216
rect 29 182 45 216
rect -91 123 -57 139
rect -91 -139 -57 -123
rect 57 123 91 139
rect 57 -139 91 -123
rect -45 -216 -29 -182
rect 29 -216 45 -182
rect -205 -284 -171 -222
rect 171 -284 205 -222
rect -205 -318 -109 -284
rect 109 -318 205 -284
<< viali >>
rect -29 182 29 216
rect -91 -123 -57 123
rect 57 -123 91 123
rect -29 -216 29 -182
<< metal1 >>
rect -41 216 41 222
rect -41 182 -29 216
rect 29 182 41 216
rect -41 176 41 182
rect -97 123 -51 135
rect -97 -123 -91 123
rect -57 -123 -51 123
rect -97 -135 -51 -123
rect 51 123 97 135
rect 51 -123 57 123
rect 91 -123 97 123
rect 51 -135 97 -123
rect -41 -182 41 -176
rect -41 -216 -29 -182
rect 29 -216 41 -182
rect -41 -222 41 -216
<< properties >>
string FIXED_BBOX -188 -301 188 301
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.35 l 0.45 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
