magic
tech sky130A
magscale 1 2
timestamp 1740547666
<< pwell >>
rect -241 -345 241 345
<< nmos >>
rect -45 -135 45 135
<< ndiff >>
rect -103 123 -45 135
rect -103 -123 -91 123
rect -57 -123 -45 123
rect -103 -135 -45 -123
rect 45 123 103 135
rect 45 -123 57 123
rect 91 -123 103 123
rect 45 -135 103 -123
<< ndiffc >>
rect -91 -123 -57 123
rect 57 -123 91 123
<< psubdiff >>
rect -205 275 -109 309
rect 109 275 205 309
rect -205 213 -171 275
rect 171 213 205 275
rect -205 -275 -171 -213
rect 171 -275 205 -213
rect -205 -309 -109 -275
rect 109 -309 205 -275
<< psubdiffcont >>
rect -109 275 109 309
rect -205 -213 -171 213
rect 171 -213 205 213
rect -109 -309 109 -275
<< poly >>
rect -45 207 45 223
rect -45 173 -29 207
rect 29 173 45 207
rect -45 135 45 173
rect -45 -173 45 -135
rect -45 -207 -29 -173
rect 29 -207 45 -173
rect -45 -223 45 -207
<< polycont >>
rect -29 173 29 207
rect -29 -207 29 -173
<< locali >>
rect -205 275 -109 309
rect 109 275 205 309
rect -205 213 -171 275
rect 171 213 205 275
rect -45 173 -29 207
rect 29 173 45 207
rect -91 123 -57 139
rect -91 -139 -57 -123
rect 57 123 91 139
rect 57 -139 91 -123
rect -45 -207 -29 -173
rect 29 -207 45 -173
rect -205 -275 -171 -213
rect 171 -275 205 -213
rect -205 -309 -109 -275
rect 109 -309 205 -275
<< viali >>
rect -29 173 29 207
rect -91 -123 -57 123
rect 57 -123 91 123
rect -29 -207 29 -173
<< metal1 >>
rect -41 207 41 213
rect -41 173 -29 207
rect 29 173 41 207
rect -41 167 41 173
rect -97 123 -51 135
rect -97 -123 -91 123
rect -57 -123 -51 123
rect -97 -135 -51 -123
rect 51 123 97 135
rect 51 -123 57 123
rect 91 -123 97 123
rect 51 -135 97 -123
rect -41 -173 41 -167
rect -41 -207 -29 -173
rect 29 -207 41 -173
rect -41 -213 41 -207
<< properties >>
string FIXED_BBOX -188 -292 188 292
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.35 l 0.450 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
